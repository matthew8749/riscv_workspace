// +FHDR--------------------------------------------------------------------------------------------------------- //
// Project ____________                                                                                           //
// File name __________ ModuleName.v                                                                              //
// Creator ____________ Yan, Wei-Ting                                                                             //
// Built Date _________ MMM-DD-YYYY                                                                               //
// Function ___________                                                                                           //
// Hierarchy __________                                                                                           //
//   Parent ___________                                                                                           //
//   Children _________                                                                                           //
// Revision history ___ Date        Author            Description                                                 //
//                  ___                                                                                           //
// -FHDR--------------------------------------------------------------------------------------------------------- //
//+...........+...................+.............................................................................. //
//3...........15..................35............................................................................. //
//`timescale 1ns/10ps

module soc_top(

  input  logic                    ref_clk_i,
  input  logic                    slow_clk_i,
  input  logic                    test_clk_i,
  input  logic                    rstn_glob_i,

);

// tag COMPONENTs and SIGNALs declaration --------------------------------------------------------------------------
  parameter                       ADR_BIT =  6;
  parameter                       DAT_BIT = 32;
  parameter                       WEN_BIT =  1;

  logic                           cen;
  logic                           wen;
  logic  [ADR_BIT-1:0]            addr;
  logic  [DAT_BIT-1:0]            din;
  logic  [DAT_BIT-1:0]            dout;


// tag OUTs assignment ---------------------------------------------------------------------------------------------
// tag INs assignment ----------------------------------------------------------------------------------------------
// tag COMBINATIONAL LOGIC -----------------------------------------------------------------------------------------
// tag COMBINATIONAL PROCESS ---------------------------------------------------------------------------------------
// tag SEQUENTIAL LOGIC --------------------------------------------------------------------------------------------
// ***********************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//                       /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *********************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

sp_ram_top i_sp_ram_top (
  .clk    ( ref_clk_i    ),
  .rst_n  ( rstn_glob_i  ),
  .CEN    ( cen          ),
  .WEN    ( wen          ),
  .addr   ( addr         ),
  .w_data ( din          ),
  .r_data ( dout         )
);

endmodule
