// +FHDR--------------------------------------------------------------------------------------------------------- //
// Project ____________                                                                                           //
// File name __________ async_fifo_SYNC_2T.sv                                                                     //
// Creator ____________ Yan, Wei-Ting                                                                             //
// Built Date _________ MMM-DD-YYYY                                                                               //
// Function ___________                                                                                           //
// Hierarchy __________                                                                                           //
//   Parent ___________                                                                                           //
//   Children _________                                                                                           //
// Revision history ___ Date        Author            Description                                                 //
//                  ___                               1.                                                          //
// -FHDR--------------------------------------------------------------------------------------------------------- //
//+...........+...................+.............................................................................. //
//3...........15..................35............................................................................. //
`timescale 1ns/10ps

module async_fifo_SYNC_2T
#(
  parameter                         SYNC_VAL_BIT = 32
)(
  input  wire                        clk,
  input  wire                        rst_n,
  input  wire [SYNC_VAL_BIT-1  : 0]  i_sync_data,
  output wire [SYNC_VAL_BIT-1  : 0]  o_sync_data
);

// tag COMPONENTs and SIGNALs declaration --------------------------------------------------------------------------
  reg   [SYNC_VAL_BIT-1 : 0]      sync_data_1t;
  reg   [SYNC_VAL_BIT-1 : 0]      sync_data_2t;

// tag OUTs assignment ---------------------------------------------------------------------------------------------
// tag OUTs assignment ---------------------------------------------------------------------------------------------
  assign  o_sync_data             = sync_data_2t;

// tag INs assignment ----------------------------------------------------------------------------------------------
// tag COMBINATIONAL LOGIC -----------------------------------------------------------------------------------------
// tag COMBINATIONAL PROCESS ---------------------------------------------------------------------------------------
// tag SEQUENTIAL LOGIC --------------------------------------------------------------------------------------------
// ***********************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//                       /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *********************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
always @ (posedge clk or negedge rst_n) begin
  if ( ~rst_n) begin
  	{sync_data_2t, sync_data_1t}  <= 'b0;
  end else begin
    {sync_data_2t, sync_data_1t}  <= {sync_data_1t, i_sync_data};


  end
end

endmodule