// This is free and unencumbered software released into the public domain.
//
// Anyone is free to copy, modify, publish, use, compile, sell, or
// distribute this software, either in source code form or as a compiled
// binary, for any purpose, commercial or non-commercial, and by any
// means.

`timescale 1 ns / 1 ps

module testbench_ez;
  reg clk = 1;
  reg resetn = 0;
  wire trap;

  always #5 clk = ~clk;

  initial begin
    $fsdbDumpfile("testbench_ez.fsdb");
    $fsdbDumpvars(0, testbench_ez, "+mda");
    $fsdbDumpMDA();
    repeat (100) @(posedge clk);
    resetn <= 1;
    repeat (100) @(posedge clk);
    $finish;
  end

  wire mem_valid;
  wire mem_instr;
  reg mem_ready;
  wire [31:0] mem_addr;
  wire [31:0] mem_wdata;
  wire [3:0] mem_wstrb;
  reg  [31:0] mem_rdata;

  always @(posedge clk) begin
    if (mem_valid && mem_ready) begin
      if (mem_instr)
        $display("ifetch 0x%08x: 0x%08x", mem_addr, mem_rdata);
      else if (mem_wstrb)
        $display("write  0x%08x: 0x%08x (wstrb=%b)", mem_addr, mem_wdata, mem_wstrb);
      else
        $display("read   0x%08x: 0x%08x", mem_addr, mem_rdata);
    end
  end

  picorv32 #(
  ) U0_picorv32 (
    .clk         (clk        ),
    .resetn      (resetn     ),
    .trap        (trap       ),
    .mem_valid   (mem_valid  ), // o
    .mem_instr   (mem_instr  ), // o
    .mem_ready   (mem_ready  ),   // i
    .mem_addr    (mem_addr   ), // o
    .mem_wdata   (mem_wdata  ), // o
    .mem_wstrb   (mem_wstrb  ), // o  //Write Strobe
    .mem_rdata   (mem_rdata  )    // i
  );

  reg [31:0] memory [0:255];

  initial begin
    memory[0] = 32'h 3fc00093; //       li      x1,1020           32'b 0011_1111_1100_ 0000_0 000_ 0000_1 001_0011        =====> addi rd, rs1, imm ;   addi x1, x0 1020
    memory[1] = 32'h 0000a023; //       sw      x0,0(x1)          32'b 0000_0000_0000_0000_1010_0000_0010_0011            =====> SW rs2, offset(rs1)
    memory[2] = 32'h 0000a103; // loop: lw      x2,0(x1)          32'b 0000_0000_0000_0000_1010_0001_0000_0011
    memory[3] = 32'h 00110113; //       addi    x2,x2,1           32'b 0000_0000_0001_0001_0000_0001_0001_0011
    memory[4] = 32'h 0020a023; //       sw      x2,0(x1)          32'b 0000_0000_0010_0000_1010_0000_0010_0011
    memory[5] = 32'h ff5ff06f; //       j       <loop>            32'b 1111_1111_0101_1111_1111_ 0000_0 110_1111            ======> jal x0, offset
  end

  always @(posedge clk) begin
    mem_ready <= 0;
    if (mem_valid && !mem_ready) begin        // "Received request" && "not yet responded ready"
      if (mem_addr < 1024) begin
        mem_ready <= 1;
        mem_rdata <= memory[mem_addr >> 2];
        if (mem_wstrb[0]) memory[mem_addr >> 2][ 7: 0] <= mem_wdata[ 7: 0];
        if (mem_wstrb[1]) memory[mem_addr >> 2][15: 8] <= mem_wdata[15: 8];
        if (mem_wstrb[2]) memory[mem_addr >> 2][23:16] <= mem_wdata[23:16];
        if (mem_wstrb[3]) memory[mem_addr >> 2][31:24] <= mem_wdata[31:24];
      end
      /* add memory-mapped IO here */
    end
  end
endmodule
