// +FHDR--------------------------------------------------------------------------------------------------------- //
// Project ____________                                                                                           //
// File name __________ sim_ram_top.sv                                                                              //
// Creator ____________ Yan, Wei-Ting                                                                             //
// Built Date _________ MMM-DD-YYYY                                                                               //
// Function ___________                                                                                           //
// Hierarchy __________                                                                                           //
//   Parent ___________                                                                                           //
//   Children _________                                                                                           //
// Revision history ___ Date        Author            Description                                                 //
//                  ___                                                                                           //
// -FHDR--------------------------------------------------------------------------------------------------------- //
//+...........+...................+.............................................................................. //
//3...........15..................35............................................................................. //
`timescale 1ns/10ps

module sp_ram_top #(
  parameter                       ADR_BIT =  6,
  parameter                       DAT_BIT = 32,
  parameter                       WEN_BIT =  1
)(
  input  logic                    clk,
  input  logic                    rst_n,
  input  logic [WEN_BIT-1: 0]     CEN,
  input  logic [WEN_BIT-1: 0]     WEN,
  input  logic [ADR_BIT-1: 0]     addr,
  input  logic [DAT_BIT-1: 0]     w_data,
  output logic [DAT_BIT-1: 0]     r_data
);

// tag COMPONENTs and SIGNALs declaration --------------------------------------------------------------------------
  logic [DAT_BIT-1: 0]            Q;
// tag OUTs assignment ---------------------------------------------------------------------------------------------
  assign      r_data            = Q;
// tag INs assignment ----------------------------------------------------------------------------------------------
// tag COMBINATIONAL LOGIC -----------------------------------------------------------------------------------------
// tag COMBINATIONAL PROCESS ---------------------------------------------------------------------------------------
// tag SEQUENTIAL LOGIC --------------------------------------------------------------------------------------------

// ***********************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//                       /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *********************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

RF1SHD_64x32 i_RF1SHD_64x32 (
  .CLK ( clk      ),
  .CEN ( CEN      ),
  .WEN ( WEN      ),
  .A   ( addr     ),
  .D   ( w_data   ),
  .Q   ( Q        )
);

endmodule