// +FHDR--------------------------------------------------------------------------------------------------------- //
// Project ____________                                                                                           //
// File name __________ linebuffer_1x640x8.sv                                                                     //
// Creator ____________ Yan, Wei-Ting                                                                             //
// Built Date _________ MMM-DD-YYYY                                                                               //
// Function ___________                                                                                           //
// Hierarchy __________                                                                                           //
//   Parent ___________                                                                                           //
//   Children _________                                                                                           //
// Revision history ___ Date        Author            Description                                                 //
//                  ___                                                                                           //
// -FHDR--------------------------------------------------------------------------------------------------------- //
//+...........+...................+.............................................................................. //
//3...........15..................35............................................................................. //
`timescale 1ns/10ps

module linebuffer_1x640x8(
  input   wire                    clk,
  input   wire                    rst_n,
  input   wire                    wr_en,
  input   wire                    rd_en,
  input   wire [ 9: 0]            addr,
  input   wire [ 7: 0]            data_in,
  output  wire [ 7: 0]            data_out
);

// tag COMPONENTs and SIGNALs declaration --------------------------------------------------------------------------
  integer                         i;

  reg  [ 7: 0]                    ram [ 639: 0];
  reg  [ 7: 0]                    bt_data_out;

// tag OUTs assignment ---------------------------------------------------------------------------------------------
  assign data_out                 = bt_data_out;

// tag INs assignment ----------------------------------------------------------------------------------------------
// tag COMBINATIONAL LOGIC -----------------------------------------------------------------------------------------
// tag COMBINATIONAL PROCESS ---------------------------------------------------------------------------------------
// tag SEQUENTIAL LOGIC --------------------------------------------------------------------------------------------
// ***********************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//                       /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *********************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****
always @ ( posedge clk or negedge rst_n ) begin
  if ( ~rst_n ) begin
    for ( i = 0; i < 10'd640; i++) begin
      ram[i] <= 8'b0;
    end
  end else begin
    ram[addr]  <= (wr_en) ? data_in  : ram[addr];


  end
end

always @ ( posedge clk or negedge rst_n ) begin
  if ( ~rst_n ) begin
    bt_data_out <= 8'b0;
  end else begin
    bt_data_out <= (rd_en) ? ram[addr] : data_in;


  end
end


endmodule



