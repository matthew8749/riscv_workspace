// +FHDR--------------------------------------------------------------------------------------------------------- //
// Project ____________                                                                                           //
// File name __________ ram_1port_mods.sv                                                                              //
// Creator ____________ Yan, Wei-Ting                                                                             //
// Built Date _________ May-19-2025                                                                               //
// Function ___________                                                                                           //
// Hierarchy __________                                                                                           //
//   Parent ___________                                                                                           //
//   Children _________                                                                                           //
// Revision history ___ Date        Author            Description                                                 //
//                  ___                                                                                           //
// -FHDR--------------------------------------------------------------------------------------------------------- //
//+...........+...................+.............................................................................. //
//3...........15..................35............................................................................. //
`timescale 1ns/1ps

module ram_1port_mod
#(
  parameter                       ADR_BIT =  4,
  parameter                       DAT_BIT = 32,
  parameter                       WEN_BIT =  1
)(
  input  wire                     clk,
  input  wire                     rst_n,
  input  wire [WEN_BIT-1: 0]      en,
  input  wire [ADR_BIT-1: 0]      addr,
  input  wire [DAT_BIT-1: 0]      w_data,
  output wire [DAT_BIT-1: 0]      r_data
);

// tag COMPONENTs and SIGNALs declaration --------------------------------------------------------------------------

// tag OUTs assignment ---------------------------------------------------------------------------------------------
// tag INs assignment ----------------------------------------------------------------------------------------------
// tag COMBINATIONAL LOGIC -----------------------------------------------------------------------------------------
// tag COMBINATIONAL PROCESS ---------------------------------------------------------------------------------------
// tag SEQUENTIAL LOGIC --------------------------------------------------------------------------------------------
// ***********************/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**\**\****/**/**
//                       /**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/****\**\**/**/***
// *********************/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/******\**\/**/****

always @ (posedge XCLK or negedge RstN) begin
  if (!RstN) begin
  end else begin

  end
end


endmodule